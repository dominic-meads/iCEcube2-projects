library ieee;
use ieee.std_logic_1164.all;

-- add file "vcomponent_vital.vhd" to modelsim project
-- found in <install_dir>\iCEcube2.2020.12\vhdl
-- compile before this entity
library work;
use work.vcomponent_vital.all; 

entity ram512x8 is
  port (
    WADDR : in std_logic_vector(8 downto 0);
    WCLK  : in std_logic;
    WCLKE : in std_logic;
    WDATA : in std_logic_vector(7 downto 0);
    WE    : in std_logic;
    RADDR : in std_logic_vector(8 downto 0);
    RCLK  : in std_logic;
    RCLKE : in std_logic;
    RE    : in std_logic;
    RDATA : out std_logic_vector(7 downto 0)
  );
end entity;

architecture rtl of ram512x8 is 

begin 

  ram512x8_inst : SB_RAM512x8 
  generic map ( 
    INIT_0 => X"0000000000000000000000000000000000000000000000000000000000000000", 
    INIT_1 => X"0000000000000000000000000000000000000000000000000000000000000000", 
    INIT_2 => X"0000000000000000000000000000000000000000000000000000000000000000", 
    INIT_3 => X"0000000000000000000000000000000000000000000000000000000000000000", 
    INIT_4 => X"0000000000000000000000000000000000000000000000000000000000000000", 
    INIT_5 => X"0000000000000000000000000000000000000000000000000000000000000000", 
    INIT_6 => X"0000000000000000000000000000000000000000000000000000000000000000", 
    INIT_7 => X"0000000000000000000000000000000000000000000000000000000000000000", 
    INIT_8 => X"0000000000000000000000000000000000000000000000000000000000000000", 
    INIT_9 => X"0000000000000000000000000000000000000000000000000000000000000000", 
    INIT_A => X"0000000000000000000000000000000000000000000000000000000000000000", 
    INIT_B => X"0000000000000000000000000000000000000000000000000000000000000000", 
    INIT_C => X"0000000000000000000000000000000000000000000000000000000000000000", 
    INIT_D => X"0000000000000000000000000000000000000000000000000000000000000000", 
    INIT_E => X"0000000000000000000000000000000000000000000000000000000000000000", 
    INIT_F => X"0000000000000000000000000000000000000000000000000000000000000000"
  ) 
  port map ( 
    RDATA => RDATA, 
    RADDR => RADDR, 
    RCLK => RCLK, 
    RCLKE => RCLKE, 
    RE => RE, 
    WADDR => WADDR, 
    WCLK=> WCLK,
    WCLKE => WCLKE, 
    WDATA => WDATA, 
    WE => WE 
  );

end architecture;
